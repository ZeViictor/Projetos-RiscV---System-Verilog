module somador ( input [7:0] a,b, output [7:0] saida)


endmodule 
